library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity cache is
generic(
	ram_size : INTEGER := 32768
);
port(
	clock : in std_logic;
	reset : in std_logic;
	
	-- Avalon interface --
	s_addr : in std_logic_vector (31 downto 0);
	s_read : in std_logic;
	s_readdata : out std_logic_vector (31 downto 0);
	s_write : in std_logic;
	s_writedata : in std_logic_vector (31 downto 0);
	s_waitrequest : out std_logic; 
    
	m_addr : out integer range 0 to ram_size-1;
	m_read : out std_logic;
	m_readdata : in std_logic_vector (7 downto 0);
	m_write : out std_logic;
	m_writedata : out std_logic_vector (7 downto 0);
	m_waitrequest : in std_logic
);
end cache;

architecture arch of cache is

type state_type is (start, r, w, r_memread, r_memwrite, r_memwait, w_memwrite);
signal state : state_type;
signal next_state : state_type;

--Address struct
--25 bits of tag
--5 bis of index
--2 bits of offset


-- Cache struct [32]
type cache_def is array (0 to 31) of std_logic_vector (154 downto 0);
signal cache2 : cache_def;
--1 bit valid  + 1 bit dirty + 25 bit tag + 128 bit data
-- 128 data + 25 tag + 1 dirty + 1 valid

begin
process (clock, reset)
begin
	if reset = '1' then
		state <= start;
	elsif (clock'event and clock = '1') then
		state <= next_state;
	end if;
end process;	

process (s_read, s_write, m_waitrequest, state)
	variable index : INTEGER;	
	variable Offset : INTEGER := 0;
	variable off : INTEGER := Offset - 1;
	variable count : INTEGER := 0;
	variable addr : std_logic_vector (14 downto 0);
begin
	index := to_integer(unsigned(s_addr(6 downto 2)));
	Offset := to_integer(unsigned(s_addr(1 downto 0))) + 1;
	off :=  Offset - 1;

	case state is
	
		when start =>
			s_waitrequest <= '1';
			if s_read = '1' then --READ
				next_state <= r;
			elsif s_write = '1' then --WRITE
				next_state <= w;
			else
				next_state <= start;
			end if;
			
		when r =>
			-- if valid and tags match
			if cache2(index)(154) = '1' and cache2(index)(152 downto 128) = s_addr (31 downto 7) then --HIT
				s_readdata <= cache2(index)(127 downto 0) ((Offset * 32) -1 downto 32*off);
				s_waitrequest <= '0';
				next_state <= start;
			elsif cache2(index)(153) = '1' then --MISS DIRTY
				next_state <= r_memwrite;
			elsif cache2(index)(153) = '0' or  cache2(index)(153) = 'U' then --MISS CLEAN
				next_state <= r_memread;
			else
				next_state <= r;
			end if;
			
		when r_memwrite =>
			if count < 4 and m_waitrequest = '1' and next_state /= r_memread then -- EVICT
				addr := cache2(index)(135 downto 128) & s_addr (6 downto 0);
				m_addr <= to_integer(unsigned (addr)) + count ;
				m_write <= '1';
				m_read <= '0';
				m_writedata <= cache2(index)(127 downto 0) ((count * 8) + 7 + 32*off downto  (count * 8) + 32*off);
				count := count + 1;
				next_state <= r_memwrite;
			elsif count = 4 then -- NOW READ FROM MEM
				count := 0;
				next_state <=r_memread;
			else
				m_write <= '0';
				next_state <= r_memwrite;
			end if;
			
		when r_memread =>
			if m_waitrequest = '1' then -- READ FROM MEM FIRST PART
				m_addr <= to_integer(unsigned(s_addr (14 downto 0))) + count;
				m_read <= '1';
				m_write <= '0';
				next_state <= r_memwait;
			else
				next_state <= r_memread;
			end if;
			
		when r_memwait =>
			if count < 3 and m_waitrequest = '0' then -- READ FROM MEM SECOND PART
				cache2(index)(127 downto 0)((count * 8) + 7 + 32*off downto  (count * 8) + 32*off) <= m_readdata;
				count := count + 1;
				m_read <= '0';
				next_state <= r_memread;
			elsif count = 3 and m_waitrequest = '0' then -- EXTRA CYCLE TO ENSURE CACHE IS READ FIRST
				cache2(index)(127 downto 0)((count * 8) + 7 + 32*off downto  (count * 8) + 32*off) <= m_readdata;
				count := count + 1;
				m_read <= '0';
				next_state <= r_memwait;
			elsif count = 4 then -- PLACE DATA READ FROM MEM ONTO OUTPUT
				s_readdata <= cache2(index)(127 downto 0) ((Offset * 32) -1 downto 32*off);
				cache2(index)(152 downto 128) <= s_addr (31 downto 7); --Tag
				cache2(index)(154) <= '1'; --Valid
				cache2(index)(153) <= '0'; --Clean
				m_read <= '0';
				m_write <= '0';
				s_waitrequest <= '0';
				count := 0;
				next_state <= start;
			else
				next_state <= r_memwait;
			end if;
		
		when w =>
			if cache2(index)(153) = '1' and next_state /= start and ( cache2(index)(154) /= '1' or cache2(index)(152 downto 128) /= s_addr (31 downto 7)) then --DIRTY AND MISS
				next_state <= w_memwrite;
			else
				cache2(index)(153) <= '1'; -- DIRTY	
				cache2(index)(154) <= '1'; --Valid
				cache2(index)(127 downto 0)((Offset * 32) -1 downto 32*off) <= s_writedata; --DATA
				cache2(index)(152 downto 128) <= s_addr (31 downto 7); --TAG
				s_waitrequest <= '0';
				next_state <= start;
					
				end if;
		
		when w_memwrite => 	
			if count < 4 and m_waitrequest = '1' then -- EVICT
				addr := cache2(index)(135 downto 128) & s_addr (6 downto 0);
				m_addr <= to_integer(unsigned (addr)) + count ;
				m_write <= '1';
				m_read <= '0';
				m_writedata <= cache2(index)(127 downto 0) ((count * 8) + 7 + 32*off downto  (count * 8) + 32*off);
				count := count + 1;
				next_state <= w_memwrite;
			elsif count = 4 then --WRITE TO CACHE AND SET CONTROL BITS
				cache2(index)(127 downto 0)((Offset * 32) -1 downto 32*off) <= s_writedata (31 downto 0); --DATA  
				cache2(index)(152 downto 128) <= s_addr (31 downto 7); --TAG
				cache2(index)(153) <= '1'; --DIRTY
				cache2(index)(154) <= '1'; --Valid
				count := 0;
				s_waitrequest <= '0';
				m_write <= '0';
				next_state <=start;
			else
				m_write <= '0';
				next_state <= w_memwrite;
			end if;
	end case;
end process;


end arch;